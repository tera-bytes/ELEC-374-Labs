library verilog;
use verilog.vl_types.all;
entity testBusMux_tb is
end testBusMux_tb;
