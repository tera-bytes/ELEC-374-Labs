library verilog;
use verilog.vl_types.all;
entity select_encode_tb is
end select_encode_tb;
