library verilog;
use verilog.vl_types.all;
entity CON_FF_tb is
end CON_FF_tb;
